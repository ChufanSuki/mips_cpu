`define PC_HASH_BITS = 3
`define PHT_INDEX_BITS = 7
